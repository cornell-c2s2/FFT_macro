magic
tech sky130A
magscale 1 2
timestamp 1682993207
<< obsli1 >>
rect 1104 2159 558808 349809
<< obsm1 >>
rect 934 76 559070 349840
<< metal2 >>
rect 8390 0 8446 800
rect 9494 0 9550 800
rect 10598 0 10654 800
rect 11702 0 11758 800
rect 12806 0 12862 800
rect 13910 0 13966 800
rect 15014 0 15070 800
rect 16118 0 16174 800
rect 17222 0 17278 800
rect 18326 0 18382 800
rect 19430 0 19486 800
rect 20534 0 20590 800
rect 21638 0 21694 800
rect 22742 0 22798 800
rect 23846 0 23902 800
rect 24950 0 25006 800
rect 26054 0 26110 800
rect 27158 0 27214 800
rect 28262 0 28318 800
rect 29366 0 29422 800
rect 30470 0 30526 800
rect 31574 0 31630 800
rect 32678 0 32734 800
rect 33782 0 33838 800
rect 34886 0 34942 800
rect 35990 0 36046 800
rect 37094 0 37150 800
rect 38198 0 38254 800
rect 39302 0 39358 800
rect 40406 0 40462 800
rect 41510 0 41566 800
rect 42614 0 42670 800
rect 43718 0 43774 800
rect 44822 0 44878 800
rect 45926 0 45982 800
rect 47030 0 47086 800
rect 48134 0 48190 800
rect 49238 0 49294 800
rect 50342 0 50398 800
rect 51446 0 51502 800
rect 52550 0 52606 800
rect 53654 0 53710 800
rect 54758 0 54814 800
rect 55862 0 55918 800
rect 56966 0 57022 800
rect 58070 0 58126 800
rect 59174 0 59230 800
rect 60278 0 60334 800
rect 61382 0 61438 800
rect 62486 0 62542 800
rect 63590 0 63646 800
rect 64694 0 64750 800
rect 65798 0 65854 800
rect 66902 0 66958 800
rect 68006 0 68062 800
rect 69110 0 69166 800
rect 70214 0 70270 800
rect 71318 0 71374 800
rect 72422 0 72478 800
rect 73526 0 73582 800
rect 74630 0 74686 800
rect 75734 0 75790 800
rect 76838 0 76894 800
rect 77942 0 77998 800
rect 79046 0 79102 800
rect 80150 0 80206 800
rect 81254 0 81310 800
rect 82358 0 82414 800
rect 83462 0 83518 800
rect 84566 0 84622 800
rect 85670 0 85726 800
rect 86774 0 86830 800
rect 87878 0 87934 800
rect 88982 0 89038 800
rect 90086 0 90142 800
rect 91190 0 91246 800
rect 92294 0 92350 800
rect 93398 0 93454 800
rect 94502 0 94558 800
rect 95606 0 95662 800
rect 96710 0 96766 800
rect 97814 0 97870 800
rect 98918 0 98974 800
rect 100022 0 100078 800
rect 101126 0 101182 800
rect 102230 0 102286 800
rect 103334 0 103390 800
rect 104438 0 104494 800
rect 105542 0 105598 800
rect 106646 0 106702 800
rect 107750 0 107806 800
rect 108854 0 108910 800
rect 109958 0 110014 800
rect 111062 0 111118 800
rect 112166 0 112222 800
rect 113270 0 113326 800
rect 114374 0 114430 800
rect 115478 0 115534 800
rect 116582 0 116638 800
rect 117686 0 117742 800
rect 118790 0 118846 800
rect 119894 0 119950 800
rect 120998 0 121054 800
rect 122102 0 122158 800
rect 123206 0 123262 800
rect 124310 0 124366 800
rect 125414 0 125470 800
rect 126518 0 126574 800
rect 127622 0 127678 800
rect 128726 0 128782 800
rect 129830 0 129886 800
rect 130934 0 130990 800
rect 132038 0 132094 800
rect 133142 0 133198 800
rect 134246 0 134302 800
rect 135350 0 135406 800
rect 136454 0 136510 800
rect 137558 0 137614 800
rect 138662 0 138718 800
rect 139766 0 139822 800
rect 140870 0 140926 800
rect 141974 0 142030 800
rect 143078 0 143134 800
rect 144182 0 144238 800
rect 145286 0 145342 800
rect 146390 0 146446 800
rect 147494 0 147550 800
rect 148598 0 148654 800
rect 149702 0 149758 800
rect 150806 0 150862 800
rect 151910 0 151966 800
rect 153014 0 153070 800
rect 154118 0 154174 800
rect 155222 0 155278 800
rect 156326 0 156382 800
rect 157430 0 157486 800
rect 158534 0 158590 800
rect 159638 0 159694 800
rect 160742 0 160798 800
rect 161846 0 161902 800
rect 162950 0 163006 800
rect 164054 0 164110 800
rect 165158 0 165214 800
rect 166262 0 166318 800
rect 167366 0 167422 800
rect 168470 0 168526 800
rect 169574 0 169630 800
rect 170678 0 170734 800
rect 171782 0 171838 800
rect 172886 0 172942 800
rect 173990 0 174046 800
rect 175094 0 175150 800
rect 176198 0 176254 800
rect 177302 0 177358 800
rect 178406 0 178462 800
rect 179510 0 179566 800
rect 180614 0 180670 800
rect 181718 0 181774 800
rect 182822 0 182878 800
rect 183926 0 183982 800
rect 185030 0 185086 800
rect 186134 0 186190 800
rect 187238 0 187294 800
rect 188342 0 188398 800
rect 189446 0 189502 800
rect 190550 0 190606 800
rect 191654 0 191710 800
rect 192758 0 192814 800
rect 193862 0 193918 800
rect 194966 0 195022 800
rect 196070 0 196126 800
rect 197174 0 197230 800
rect 198278 0 198334 800
rect 199382 0 199438 800
rect 200486 0 200542 800
rect 201590 0 201646 800
rect 202694 0 202750 800
rect 203798 0 203854 800
rect 204902 0 204958 800
rect 206006 0 206062 800
rect 207110 0 207166 800
rect 208214 0 208270 800
rect 209318 0 209374 800
rect 210422 0 210478 800
rect 211526 0 211582 800
rect 212630 0 212686 800
rect 213734 0 213790 800
rect 214838 0 214894 800
rect 215942 0 215998 800
rect 217046 0 217102 800
rect 218150 0 218206 800
rect 219254 0 219310 800
rect 220358 0 220414 800
rect 221462 0 221518 800
rect 222566 0 222622 800
rect 223670 0 223726 800
rect 224774 0 224830 800
rect 225878 0 225934 800
rect 226982 0 227038 800
rect 228086 0 228142 800
rect 229190 0 229246 800
rect 230294 0 230350 800
rect 231398 0 231454 800
rect 232502 0 232558 800
rect 233606 0 233662 800
rect 234710 0 234766 800
rect 235814 0 235870 800
rect 236918 0 236974 800
rect 238022 0 238078 800
rect 239126 0 239182 800
rect 240230 0 240286 800
rect 241334 0 241390 800
rect 242438 0 242494 800
rect 243542 0 243598 800
rect 244646 0 244702 800
rect 245750 0 245806 800
rect 246854 0 246910 800
rect 247958 0 248014 800
rect 249062 0 249118 800
rect 250166 0 250222 800
rect 251270 0 251326 800
rect 252374 0 252430 800
rect 253478 0 253534 800
rect 254582 0 254638 800
rect 255686 0 255742 800
rect 256790 0 256846 800
rect 257894 0 257950 800
rect 258998 0 259054 800
rect 260102 0 260158 800
rect 261206 0 261262 800
rect 262310 0 262366 800
rect 263414 0 263470 800
rect 264518 0 264574 800
rect 265622 0 265678 800
rect 266726 0 266782 800
rect 267830 0 267886 800
rect 268934 0 268990 800
rect 270038 0 270094 800
rect 271142 0 271198 800
rect 272246 0 272302 800
rect 273350 0 273406 800
rect 274454 0 274510 800
rect 275558 0 275614 800
rect 276662 0 276718 800
rect 277766 0 277822 800
rect 278870 0 278926 800
rect 279974 0 280030 800
rect 281078 0 281134 800
rect 282182 0 282238 800
rect 283286 0 283342 800
rect 284390 0 284446 800
rect 285494 0 285550 800
rect 286598 0 286654 800
rect 287702 0 287758 800
rect 288806 0 288862 800
rect 289910 0 289966 800
rect 291014 0 291070 800
rect 292118 0 292174 800
rect 293222 0 293278 800
rect 294326 0 294382 800
rect 295430 0 295486 800
rect 296534 0 296590 800
rect 297638 0 297694 800
rect 298742 0 298798 800
rect 299846 0 299902 800
rect 300950 0 301006 800
rect 302054 0 302110 800
rect 303158 0 303214 800
rect 304262 0 304318 800
rect 305366 0 305422 800
rect 306470 0 306526 800
rect 307574 0 307630 800
rect 308678 0 308734 800
rect 309782 0 309838 800
rect 310886 0 310942 800
rect 311990 0 312046 800
rect 313094 0 313150 800
rect 314198 0 314254 800
rect 315302 0 315358 800
rect 316406 0 316462 800
rect 317510 0 317566 800
rect 318614 0 318670 800
rect 319718 0 319774 800
rect 320822 0 320878 800
rect 321926 0 321982 800
rect 323030 0 323086 800
rect 324134 0 324190 800
rect 325238 0 325294 800
rect 326342 0 326398 800
rect 327446 0 327502 800
rect 328550 0 328606 800
rect 329654 0 329710 800
rect 330758 0 330814 800
rect 331862 0 331918 800
rect 332966 0 333022 800
rect 334070 0 334126 800
rect 335174 0 335230 800
rect 336278 0 336334 800
rect 337382 0 337438 800
rect 338486 0 338542 800
rect 339590 0 339646 800
rect 340694 0 340750 800
rect 341798 0 341854 800
rect 342902 0 342958 800
rect 344006 0 344062 800
rect 345110 0 345166 800
rect 346214 0 346270 800
rect 347318 0 347374 800
rect 348422 0 348478 800
rect 349526 0 349582 800
rect 350630 0 350686 800
rect 351734 0 351790 800
rect 352838 0 352894 800
rect 353942 0 353998 800
rect 355046 0 355102 800
rect 356150 0 356206 800
rect 357254 0 357310 800
rect 358358 0 358414 800
rect 359462 0 359518 800
rect 360566 0 360622 800
rect 361670 0 361726 800
rect 362774 0 362830 800
rect 363878 0 363934 800
rect 364982 0 365038 800
rect 366086 0 366142 800
rect 367190 0 367246 800
rect 368294 0 368350 800
rect 369398 0 369454 800
rect 370502 0 370558 800
rect 371606 0 371662 800
rect 372710 0 372766 800
rect 373814 0 373870 800
rect 374918 0 374974 800
rect 376022 0 376078 800
rect 377126 0 377182 800
rect 378230 0 378286 800
rect 379334 0 379390 800
rect 380438 0 380494 800
rect 381542 0 381598 800
rect 382646 0 382702 800
rect 383750 0 383806 800
rect 384854 0 384910 800
rect 385958 0 386014 800
rect 387062 0 387118 800
rect 388166 0 388222 800
rect 389270 0 389326 800
rect 390374 0 390430 800
rect 391478 0 391534 800
rect 392582 0 392638 800
rect 393686 0 393742 800
rect 394790 0 394846 800
rect 395894 0 395950 800
rect 396998 0 397054 800
rect 398102 0 398158 800
rect 399206 0 399262 800
rect 400310 0 400366 800
rect 401414 0 401470 800
rect 402518 0 402574 800
rect 403622 0 403678 800
rect 404726 0 404782 800
rect 405830 0 405886 800
rect 406934 0 406990 800
rect 408038 0 408094 800
rect 409142 0 409198 800
rect 410246 0 410302 800
rect 411350 0 411406 800
rect 412454 0 412510 800
rect 413558 0 413614 800
rect 414662 0 414718 800
rect 415766 0 415822 800
rect 416870 0 416926 800
rect 417974 0 418030 800
rect 419078 0 419134 800
rect 420182 0 420238 800
rect 421286 0 421342 800
rect 422390 0 422446 800
rect 423494 0 423550 800
rect 424598 0 424654 800
rect 425702 0 425758 800
rect 426806 0 426862 800
rect 427910 0 427966 800
rect 429014 0 429070 800
rect 430118 0 430174 800
rect 431222 0 431278 800
rect 432326 0 432382 800
rect 433430 0 433486 800
rect 434534 0 434590 800
rect 435638 0 435694 800
rect 436742 0 436798 800
rect 437846 0 437902 800
rect 438950 0 439006 800
rect 440054 0 440110 800
rect 441158 0 441214 800
rect 442262 0 442318 800
rect 443366 0 443422 800
rect 444470 0 444526 800
rect 445574 0 445630 800
rect 446678 0 446734 800
rect 447782 0 447838 800
rect 448886 0 448942 800
rect 449990 0 450046 800
rect 451094 0 451150 800
rect 452198 0 452254 800
rect 453302 0 453358 800
rect 454406 0 454462 800
rect 455510 0 455566 800
rect 456614 0 456670 800
rect 457718 0 457774 800
rect 458822 0 458878 800
rect 459926 0 459982 800
rect 461030 0 461086 800
rect 462134 0 462190 800
rect 463238 0 463294 800
rect 464342 0 464398 800
rect 465446 0 465502 800
rect 466550 0 466606 800
rect 467654 0 467710 800
rect 468758 0 468814 800
rect 469862 0 469918 800
rect 470966 0 471022 800
rect 472070 0 472126 800
rect 473174 0 473230 800
rect 474278 0 474334 800
rect 475382 0 475438 800
rect 476486 0 476542 800
rect 477590 0 477646 800
rect 478694 0 478750 800
rect 479798 0 479854 800
rect 480902 0 480958 800
rect 482006 0 482062 800
rect 483110 0 483166 800
rect 484214 0 484270 800
rect 485318 0 485374 800
rect 486422 0 486478 800
rect 487526 0 487582 800
rect 488630 0 488686 800
rect 489734 0 489790 800
rect 490838 0 490894 800
rect 491942 0 491998 800
rect 493046 0 493102 800
rect 494150 0 494206 800
rect 495254 0 495310 800
rect 496358 0 496414 800
rect 497462 0 497518 800
rect 498566 0 498622 800
rect 499670 0 499726 800
rect 500774 0 500830 800
rect 501878 0 501934 800
rect 502982 0 503038 800
rect 504086 0 504142 800
rect 505190 0 505246 800
rect 506294 0 506350 800
rect 507398 0 507454 800
rect 508502 0 508558 800
rect 509606 0 509662 800
rect 510710 0 510766 800
rect 511814 0 511870 800
rect 512918 0 512974 800
rect 514022 0 514078 800
rect 515126 0 515182 800
rect 516230 0 516286 800
rect 517334 0 517390 800
rect 518438 0 518494 800
rect 519542 0 519598 800
rect 520646 0 520702 800
rect 521750 0 521806 800
rect 522854 0 522910 800
rect 523958 0 524014 800
rect 525062 0 525118 800
rect 526166 0 526222 800
rect 527270 0 527326 800
rect 528374 0 528430 800
rect 529478 0 529534 800
rect 530582 0 530638 800
rect 531686 0 531742 800
rect 532790 0 532846 800
rect 533894 0 533950 800
rect 534998 0 535054 800
rect 536102 0 536158 800
rect 537206 0 537262 800
rect 538310 0 538366 800
rect 539414 0 539470 800
rect 540518 0 540574 800
rect 541622 0 541678 800
rect 542726 0 542782 800
rect 543830 0 543886 800
rect 544934 0 544990 800
rect 546038 0 546094 800
rect 547142 0 547198 800
rect 548246 0 548302 800
rect 549350 0 549406 800
rect 550454 0 550510 800
rect 551558 0 551614 800
<< obsm2 >>
rect 938 856 559066 349829
rect 938 31 8334 856
rect 8502 31 9438 856
rect 9606 31 10542 856
rect 10710 31 11646 856
rect 11814 31 12750 856
rect 12918 31 13854 856
rect 14022 31 14958 856
rect 15126 31 16062 856
rect 16230 31 17166 856
rect 17334 31 18270 856
rect 18438 31 19374 856
rect 19542 31 20478 856
rect 20646 31 21582 856
rect 21750 31 22686 856
rect 22854 31 23790 856
rect 23958 31 24894 856
rect 25062 31 25998 856
rect 26166 31 27102 856
rect 27270 31 28206 856
rect 28374 31 29310 856
rect 29478 31 30414 856
rect 30582 31 31518 856
rect 31686 31 32622 856
rect 32790 31 33726 856
rect 33894 31 34830 856
rect 34998 31 35934 856
rect 36102 31 37038 856
rect 37206 31 38142 856
rect 38310 31 39246 856
rect 39414 31 40350 856
rect 40518 31 41454 856
rect 41622 31 42558 856
rect 42726 31 43662 856
rect 43830 31 44766 856
rect 44934 31 45870 856
rect 46038 31 46974 856
rect 47142 31 48078 856
rect 48246 31 49182 856
rect 49350 31 50286 856
rect 50454 31 51390 856
rect 51558 31 52494 856
rect 52662 31 53598 856
rect 53766 31 54702 856
rect 54870 31 55806 856
rect 55974 31 56910 856
rect 57078 31 58014 856
rect 58182 31 59118 856
rect 59286 31 60222 856
rect 60390 31 61326 856
rect 61494 31 62430 856
rect 62598 31 63534 856
rect 63702 31 64638 856
rect 64806 31 65742 856
rect 65910 31 66846 856
rect 67014 31 67950 856
rect 68118 31 69054 856
rect 69222 31 70158 856
rect 70326 31 71262 856
rect 71430 31 72366 856
rect 72534 31 73470 856
rect 73638 31 74574 856
rect 74742 31 75678 856
rect 75846 31 76782 856
rect 76950 31 77886 856
rect 78054 31 78990 856
rect 79158 31 80094 856
rect 80262 31 81198 856
rect 81366 31 82302 856
rect 82470 31 83406 856
rect 83574 31 84510 856
rect 84678 31 85614 856
rect 85782 31 86718 856
rect 86886 31 87822 856
rect 87990 31 88926 856
rect 89094 31 90030 856
rect 90198 31 91134 856
rect 91302 31 92238 856
rect 92406 31 93342 856
rect 93510 31 94446 856
rect 94614 31 95550 856
rect 95718 31 96654 856
rect 96822 31 97758 856
rect 97926 31 98862 856
rect 99030 31 99966 856
rect 100134 31 101070 856
rect 101238 31 102174 856
rect 102342 31 103278 856
rect 103446 31 104382 856
rect 104550 31 105486 856
rect 105654 31 106590 856
rect 106758 31 107694 856
rect 107862 31 108798 856
rect 108966 31 109902 856
rect 110070 31 111006 856
rect 111174 31 112110 856
rect 112278 31 113214 856
rect 113382 31 114318 856
rect 114486 31 115422 856
rect 115590 31 116526 856
rect 116694 31 117630 856
rect 117798 31 118734 856
rect 118902 31 119838 856
rect 120006 31 120942 856
rect 121110 31 122046 856
rect 122214 31 123150 856
rect 123318 31 124254 856
rect 124422 31 125358 856
rect 125526 31 126462 856
rect 126630 31 127566 856
rect 127734 31 128670 856
rect 128838 31 129774 856
rect 129942 31 130878 856
rect 131046 31 131982 856
rect 132150 31 133086 856
rect 133254 31 134190 856
rect 134358 31 135294 856
rect 135462 31 136398 856
rect 136566 31 137502 856
rect 137670 31 138606 856
rect 138774 31 139710 856
rect 139878 31 140814 856
rect 140982 31 141918 856
rect 142086 31 143022 856
rect 143190 31 144126 856
rect 144294 31 145230 856
rect 145398 31 146334 856
rect 146502 31 147438 856
rect 147606 31 148542 856
rect 148710 31 149646 856
rect 149814 31 150750 856
rect 150918 31 151854 856
rect 152022 31 152958 856
rect 153126 31 154062 856
rect 154230 31 155166 856
rect 155334 31 156270 856
rect 156438 31 157374 856
rect 157542 31 158478 856
rect 158646 31 159582 856
rect 159750 31 160686 856
rect 160854 31 161790 856
rect 161958 31 162894 856
rect 163062 31 163998 856
rect 164166 31 165102 856
rect 165270 31 166206 856
rect 166374 31 167310 856
rect 167478 31 168414 856
rect 168582 31 169518 856
rect 169686 31 170622 856
rect 170790 31 171726 856
rect 171894 31 172830 856
rect 172998 31 173934 856
rect 174102 31 175038 856
rect 175206 31 176142 856
rect 176310 31 177246 856
rect 177414 31 178350 856
rect 178518 31 179454 856
rect 179622 31 180558 856
rect 180726 31 181662 856
rect 181830 31 182766 856
rect 182934 31 183870 856
rect 184038 31 184974 856
rect 185142 31 186078 856
rect 186246 31 187182 856
rect 187350 31 188286 856
rect 188454 31 189390 856
rect 189558 31 190494 856
rect 190662 31 191598 856
rect 191766 31 192702 856
rect 192870 31 193806 856
rect 193974 31 194910 856
rect 195078 31 196014 856
rect 196182 31 197118 856
rect 197286 31 198222 856
rect 198390 31 199326 856
rect 199494 31 200430 856
rect 200598 31 201534 856
rect 201702 31 202638 856
rect 202806 31 203742 856
rect 203910 31 204846 856
rect 205014 31 205950 856
rect 206118 31 207054 856
rect 207222 31 208158 856
rect 208326 31 209262 856
rect 209430 31 210366 856
rect 210534 31 211470 856
rect 211638 31 212574 856
rect 212742 31 213678 856
rect 213846 31 214782 856
rect 214950 31 215886 856
rect 216054 31 216990 856
rect 217158 31 218094 856
rect 218262 31 219198 856
rect 219366 31 220302 856
rect 220470 31 221406 856
rect 221574 31 222510 856
rect 222678 31 223614 856
rect 223782 31 224718 856
rect 224886 31 225822 856
rect 225990 31 226926 856
rect 227094 31 228030 856
rect 228198 31 229134 856
rect 229302 31 230238 856
rect 230406 31 231342 856
rect 231510 31 232446 856
rect 232614 31 233550 856
rect 233718 31 234654 856
rect 234822 31 235758 856
rect 235926 31 236862 856
rect 237030 31 237966 856
rect 238134 31 239070 856
rect 239238 31 240174 856
rect 240342 31 241278 856
rect 241446 31 242382 856
rect 242550 31 243486 856
rect 243654 31 244590 856
rect 244758 31 245694 856
rect 245862 31 246798 856
rect 246966 31 247902 856
rect 248070 31 249006 856
rect 249174 31 250110 856
rect 250278 31 251214 856
rect 251382 31 252318 856
rect 252486 31 253422 856
rect 253590 31 254526 856
rect 254694 31 255630 856
rect 255798 31 256734 856
rect 256902 31 257838 856
rect 258006 31 258942 856
rect 259110 31 260046 856
rect 260214 31 261150 856
rect 261318 31 262254 856
rect 262422 31 263358 856
rect 263526 31 264462 856
rect 264630 31 265566 856
rect 265734 31 266670 856
rect 266838 31 267774 856
rect 267942 31 268878 856
rect 269046 31 269982 856
rect 270150 31 271086 856
rect 271254 31 272190 856
rect 272358 31 273294 856
rect 273462 31 274398 856
rect 274566 31 275502 856
rect 275670 31 276606 856
rect 276774 31 277710 856
rect 277878 31 278814 856
rect 278982 31 279918 856
rect 280086 31 281022 856
rect 281190 31 282126 856
rect 282294 31 283230 856
rect 283398 31 284334 856
rect 284502 31 285438 856
rect 285606 31 286542 856
rect 286710 31 287646 856
rect 287814 31 288750 856
rect 288918 31 289854 856
rect 290022 31 290958 856
rect 291126 31 292062 856
rect 292230 31 293166 856
rect 293334 31 294270 856
rect 294438 31 295374 856
rect 295542 31 296478 856
rect 296646 31 297582 856
rect 297750 31 298686 856
rect 298854 31 299790 856
rect 299958 31 300894 856
rect 301062 31 301998 856
rect 302166 31 303102 856
rect 303270 31 304206 856
rect 304374 31 305310 856
rect 305478 31 306414 856
rect 306582 31 307518 856
rect 307686 31 308622 856
rect 308790 31 309726 856
rect 309894 31 310830 856
rect 310998 31 311934 856
rect 312102 31 313038 856
rect 313206 31 314142 856
rect 314310 31 315246 856
rect 315414 31 316350 856
rect 316518 31 317454 856
rect 317622 31 318558 856
rect 318726 31 319662 856
rect 319830 31 320766 856
rect 320934 31 321870 856
rect 322038 31 322974 856
rect 323142 31 324078 856
rect 324246 31 325182 856
rect 325350 31 326286 856
rect 326454 31 327390 856
rect 327558 31 328494 856
rect 328662 31 329598 856
rect 329766 31 330702 856
rect 330870 31 331806 856
rect 331974 31 332910 856
rect 333078 31 334014 856
rect 334182 31 335118 856
rect 335286 31 336222 856
rect 336390 31 337326 856
rect 337494 31 338430 856
rect 338598 31 339534 856
rect 339702 31 340638 856
rect 340806 31 341742 856
rect 341910 31 342846 856
rect 343014 31 343950 856
rect 344118 31 345054 856
rect 345222 31 346158 856
rect 346326 31 347262 856
rect 347430 31 348366 856
rect 348534 31 349470 856
rect 349638 31 350574 856
rect 350742 31 351678 856
rect 351846 31 352782 856
rect 352950 31 353886 856
rect 354054 31 354990 856
rect 355158 31 356094 856
rect 356262 31 357198 856
rect 357366 31 358302 856
rect 358470 31 359406 856
rect 359574 31 360510 856
rect 360678 31 361614 856
rect 361782 31 362718 856
rect 362886 31 363822 856
rect 363990 31 364926 856
rect 365094 31 366030 856
rect 366198 31 367134 856
rect 367302 31 368238 856
rect 368406 31 369342 856
rect 369510 31 370446 856
rect 370614 31 371550 856
rect 371718 31 372654 856
rect 372822 31 373758 856
rect 373926 31 374862 856
rect 375030 31 375966 856
rect 376134 31 377070 856
rect 377238 31 378174 856
rect 378342 31 379278 856
rect 379446 31 380382 856
rect 380550 31 381486 856
rect 381654 31 382590 856
rect 382758 31 383694 856
rect 383862 31 384798 856
rect 384966 31 385902 856
rect 386070 31 387006 856
rect 387174 31 388110 856
rect 388278 31 389214 856
rect 389382 31 390318 856
rect 390486 31 391422 856
rect 391590 31 392526 856
rect 392694 31 393630 856
rect 393798 31 394734 856
rect 394902 31 395838 856
rect 396006 31 396942 856
rect 397110 31 398046 856
rect 398214 31 399150 856
rect 399318 31 400254 856
rect 400422 31 401358 856
rect 401526 31 402462 856
rect 402630 31 403566 856
rect 403734 31 404670 856
rect 404838 31 405774 856
rect 405942 31 406878 856
rect 407046 31 407982 856
rect 408150 31 409086 856
rect 409254 31 410190 856
rect 410358 31 411294 856
rect 411462 31 412398 856
rect 412566 31 413502 856
rect 413670 31 414606 856
rect 414774 31 415710 856
rect 415878 31 416814 856
rect 416982 31 417918 856
rect 418086 31 419022 856
rect 419190 31 420126 856
rect 420294 31 421230 856
rect 421398 31 422334 856
rect 422502 31 423438 856
rect 423606 31 424542 856
rect 424710 31 425646 856
rect 425814 31 426750 856
rect 426918 31 427854 856
rect 428022 31 428958 856
rect 429126 31 430062 856
rect 430230 31 431166 856
rect 431334 31 432270 856
rect 432438 31 433374 856
rect 433542 31 434478 856
rect 434646 31 435582 856
rect 435750 31 436686 856
rect 436854 31 437790 856
rect 437958 31 438894 856
rect 439062 31 439998 856
rect 440166 31 441102 856
rect 441270 31 442206 856
rect 442374 31 443310 856
rect 443478 31 444414 856
rect 444582 31 445518 856
rect 445686 31 446622 856
rect 446790 31 447726 856
rect 447894 31 448830 856
rect 448998 31 449934 856
rect 450102 31 451038 856
rect 451206 31 452142 856
rect 452310 31 453246 856
rect 453414 31 454350 856
rect 454518 31 455454 856
rect 455622 31 456558 856
rect 456726 31 457662 856
rect 457830 31 458766 856
rect 458934 31 459870 856
rect 460038 31 460974 856
rect 461142 31 462078 856
rect 462246 31 463182 856
rect 463350 31 464286 856
rect 464454 31 465390 856
rect 465558 31 466494 856
rect 466662 31 467598 856
rect 467766 31 468702 856
rect 468870 31 469806 856
rect 469974 31 470910 856
rect 471078 31 472014 856
rect 472182 31 473118 856
rect 473286 31 474222 856
rect 474390 31 475326 856
rect 475494 31 476430 856
rect 476598 31 477534 856
rect 477702 31 478638 856
rect 478806 31 479742 856
rect 479910 31 480846 856
rect 481014 31 481950 856
rect 482118 31 483054 856
rect 483222 31 484158 856
rect 484326 31 485262 856
rect 485430 31 486366 856
rect 486534 31 487470 856
rect 487638 31 488574 856
rect 488742 31 489678 856
rect 489846 31 490782 856
rect 490950 31 491886 856
rect 492054 31 492990 856
rect 493158 31 494094 856
rect 494262 31 495198 856
rect 495366 31 496302 856
rect 496470 31 497406 856
rect 497574 31 498510 856
rect 498678 31 499614 856
rect 499782 31 500718 856
rect 500886 31 501822 856
rect 501990 31 502926 856
rect 503094 31 504030 856
rect 504198 31 505134 856
rect 505302 31 506238 856
rect 506406 31 507342 856
rect 507510 31 508446 856
rect 508614 31 509550 856
rect 509718 31 510654 856
rect 510822 31 511758 856
rect 511926 31 512862 856
rect 513030 31 513966 856
rect 514134 31 515070 856
rect 515238 31 516174 856
rect 516342 31 517278 856
rect 517446 31 518382 856
rect 518550 31 519486 856
rect 519654 31 520590 856
rect 520758 31 521694 856
rect 521862 31 522798 856
rect 522966 31 523902 856
rect 524070 31 525006 856
rect 525174 31 526110 856
rect 526278 31 527214 856
rect 527382 31 528318 856
rect 528486 31 529422 856
rect 529590 31 530526 856
rect 530694 31 531630 856
rect 531798 31 532734 856
rect 532902 31 533838 856
rect 534006 31 534942 856
rect 535110 31 536046 856
rect 536214 31 537150 856
rect 537318 31 538254 856
rect 538422 31 539358 856
rect 539526 31 540462 856
rect 540630 31 541566 856
rect 541734 31 542670 856
rect 542838 31 543774 856
rect 543942 31 544878 856
rect 545046 31 545982 856
rect 546150 31 547086 856
rect 547254 31 548190 856
rect 548358 31 549294 856
rect 549462 31 550398 856
rect 550566 31 551502 856
rect 551670 31 559066 856
<< metal3 >>
rect 0 343272 800 343392
rect 559200 343272 560000 343392
rect 0 328720 800 328840
rect 559200 328720 560000 328840
rect 0 314168 800 314288
rect 559200 314168 560000 314288
rect 0 299616 800 299736
rect 559200 299616 560000 299736
rect 0 285064 800 285184
rect 559200 285064 560000 285184
rect 0 270512 800 270632
rect 559200 270512 560000 270632
rect 0 255960 800 256080
rect 559200 255960 560000 256080
rect 0 241408 800 241528
rect 559200 241408 560000 241528
rect 0 226856 800 226976
rect 559200 226856 560000 226976
rect 0 212304 800 212424
rect 559200 212304 560000 212424
rect 0 197752 800 197872
rect 559200 197752 560000 197872
rect 0 183200 800 183320
rect 559200 183200 560000 183320
rect 0 168648 800 168768
rect 559200 168648 560000 168768
rect 0 154096 800 154216
rect 559200 154096 560000 154216
rect 0 139544 800 139664
rect 559200 139544 560000 139664
rect 0 124992 800 125112
rect 559200 124992 560000 125112
rect 0 110440 800 110560
rect 559200 110440 560000 110560
rect 0 95888 800 96008
rect 559200 95888 560000 96008
rect 0 81336 800 81456
rect 559200 81336 560000 81456
rect 0 66784 800 66904
rect 559200 66784 560000 66904
rect 0 52232 800 52352
rect 559200 52232 560000 52352
rect 0 37680 800 37800
rect 559200 37680 560000 37800
rect 0 23128 800 23248
rect 559200 23128 560000 23248
rect 0 8576 800 8696
rect 559200 8576 560000 8696
<< obsm3 >>
rect 800 343472 559200 349825
rect 880 343192 559120 343472
rect 800 328920 559200 343192
rect 880 328640 559120 328920
rect 800 314368 559200 328640
rect 880 314088 559120 314368
rect 800 299816 559200 314088
rect 880 299536 559120 299816
rect 800 285264 559200 299536
rect 880 284984 559120 285264
rect 800 270712 559200 284984
rect 880 270432 559120 270712
rect 800 256160 559200 270432
rect 880 255880 559120 256160
rect 800 241608 559200 255880
rect 880 241328 559120 241608
rect 800 227056 559200 241328
rect 880 226776 559120 227056
rect 800 212504 559200 226776
rect 880 212224 559120 212504
rect 800 197952 559200 212224
rect 880 197672 559120 197952
rect 800 183400 559200 197672
rect 880 183120 559120 183400
rect 800 168848 559200 183120
rect 880 168568 559120 168848
rect 800 154296 559200 168568
rect 880 154016 559120 154296
rect 800 139744 559200 154016
rect 880 139464 559120 139744
rect 800 125192 559200 139464
rect 880 124912 559120 125192
rect 800 110640 559200 124912
rect 880 110360 559120 110640
rect 800 96088 559200 110360
rect 880 95808 559120 96088
rect 800 81536 559200 95808
rect 880 81256 559120 81536
rect 800 66984 559200 81256
rect 880 66704 559120 66984
rect 800 52432 559200 66704
rect 880 52152 559120 52432
rect 800 37880 559200 52152
rect 880 37600 559120 37880
rect 800 23328 559200 37600
rect 880 23048 559120 23328
rect 800 8776 559200 23048
rect 880 8496 559120 8776
rect 800 35 559200 8496
<< metal4 >>
rect 4208 2128 4528 349840
rect 19568 2128 19888 349840
rect 34928 2128 35248 349840
rect 50288 2128 50608 349840
rect 65648 2128 65968 349840
rect 81008 2128 81328 349840
rect 96368 2128 96688 349840
rect 111728 2128 112048 349840
rect 127088 2128 127408 349840
rect 142448 2128 142768 349840
rect 157808 2128 158128 349840
rect 173168 2128 173488 349840
rect 188528 2128 188848 349840
rect 203888 2128 204208 349840
rect 219248 2128 219568 349840
rect 234608 2128 234928 349840
rect 249968 2128 250288 349840
rect 265328 2128 265648 349840
rect 280688 2128 281008 349840
rect 296048 2128 296368 349840
rect 311408 2128 311728 349840
rect 326768 2128 327088 349840
rect 342128 2128 342448 349840
rect 357488 2128 357808 349840
rect 372848 2128 373168 349840
rect 388208 2128 388528 349840
rect 403568 2128 403888 349840
rect 418928 2128 419248 349840
rect 434288 2128 434608 349840
rect 449648 2128 449968 349840
rect 465008 2128 465328 349840
rect 480368 2128 480688 349840
rect 495728 2128 496048 349840
rect 511088 2128 511408 349840
rect 526448 2128 526768 349840
rect 541808 2128 542128 349840
rect 557168 2128 557488 349840
<< obsm4 >>
rect 230059 3163 234528 22133
rect 235008 3163 243925 22133
<< labels >>
rlabel metal3 s 559200 8576 560000 8696 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 0 255960 800 256080 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 0 212304 800 212424 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 0 168648 800 168768 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 0 124992 800 125112 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 0 81336 800 81456 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 0 37680 800 37800 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 559200 52232 560000 52352 6 io_in[1]
port 8 nsew signal input
rlabel metal3 s 559200 95888 560000 96008 6 io_in[2]
port 9 nsew signal input
rlabel metal3 s 559200 139544 560000 139664 6 io_in[3]
port 10 nsew signal input
rlabel metal3 s 559200 183200 560000 183320 6 io_in[4]
port 11 nsew signal input
rlabel metal3 s 559200 226856 560000 226976 6 io_in[5]
port 12 nsew signal input
rlabel metal3 s 559200 270512 560000 270632 6 io_in[6]
port 13 nsew signal input
rlabel metal3 s 559200 314168 560000 314288 6 io_in[7]
port 14 nsew signal input
rlabel metal3 s 0 343272 800 343392 6 io_in[8]
port 15 nsew signal input
rlabel metal3 s 0 299616 800 299736 6 io_in[9]
port 16 nsew signal input
rlabel metal3 s 559200 37680 560000 37800 6 io_oeb[0]
port 17 nsew signal output
rlabel metal3 s 0 226856 800 226976 6 io_oeb[10]
port 18 nsew signal output
rlabel metal3 s 0 183200 800 183320 6 io_oeb[11]
port 19 nsew signal output
rlabel metal3 s 0 139544 800 139664 6 io_oeb[12]
port 20 nsew signal output
rlabel metal3 s 0 95888 800 96008 6 io_oeb[13]
port 21 nsew signal output
rlabel metal3 s 0 52232 800 52352 6 io_oeb[14]
port 22 nsew signal output
rlabel metal3 s 0 8576 800 8696 6 io_oeb[15]
port 23 nsew signal output
rlabel metal3 s 559200 81336 560000 81456 6 io_oeb[1]
port 24 nsew signal output
rlabel metal3 s 559200 124992 560000 125112 6 io_oeb[2]
port 25 nsew signal output
rlabel metal3 s 559200 168648 560000 168768 6 io_oeb[3]
port 26 nsew signal output
rlabel metal3 s 559200 212304 560000 212424 6 io_oeb[4]
port 27 nsew signal output
rlabel metal3 s 559200 255960 560000 256080 6 io_oeb[5]
port 28 nsew signal output
rlabel metal3 s 559200 299616 560000 299736 6 io_oeb[6]
port 29 nsew signal output
rlabel metal3 s 559200 343272 560000 343392 6 io_oeb[7]
port 30 nsew signal output
rlabel metal3 s 0 314168 800 314288 6 io_oeb[8]
port 31 nsew signal output
rlabel metal3 s 0 270512 800 270632 6 io_oeb[9]
port 32 nsew signal output
rlabel metal3 s 559200 23128 560000 23248 6 io_out[0]
port 33 nsew signal output
rlabel metal3 s 0 241408 800 241528 6 io_out[10]
port 34 nsew signal output
rlabel metal3 s 0 197752 800 197872 6 io_out[11]
port 35 nsew signal output
rlabel metal3 s 0 154096 800 154216 6 io_out[12]
port 36 nsew signal output
rlabel metal3 s 0 110440 800 110560 6 io_out[13]
port 37 nsew signal output
rlabel metal3 s 0 66784 800 66904 6 io_out[14]
port 38 nsew signal output
rlabel metal3 s 0 23128 800 23248 6 io_out[15]
port 39 nsew signal output
rlabel metal3 s 559200 66784 560000 66904 6 io_out[1]
port 40 nsew signal output
rlabel metal3 s 559200 110440 560000 110560 6 io_out[2]
port 41 nsew signal output
rlabel metal3 s 559200 154096 560000 154216 6 io_out[3]
port 42 nsew signal output
rlabel metal3 s 559200 197752 560000 197872 6 io_out[4]
port 43 nsew signal output
rlabel metal3 s 559200 241408 560000 241528 6 io_out[5]
port 44 nsew signal output
rlabel metal3 s 559200 285064 560000 285184 6 io_out[6]
port 45 nsew signal output
rlabel metal3 s 559200 328720 560000 328840 6 io_out[7]
port 46 nsew signal output
rlabel metal3 s 0 328720 800 328840 6 io_out[8]
port 47 nsew signal output
rlabel metal3 s 0 285064 800 285184 6 io_out[9]
port 48 nsew signal output
rlabel metal2 s 549350 0 549406 800 6 irq[0]
port 49 nsew signal output
rlabel metal2 s 550454 0 550510 800 6 irq[1]
port 50 nsew signal output
rlabel metal2 s 551558 0 551614 800 6 irq[2]
port 51 nsew signal output
rlabel metal2 s 125414 0 125470 800 6 la_data_in[0]
port 52 nsew signal input
rlabel metal2 s 456614 0 456670 800 6 la_data_in[100]
port 53 nsew signal input
rlabel metal2 s 459926 0 459982 800 6 la_data_in[101]
port 54 nsew signal input
rlabel metal2 s 463238 0 463294 800 6 la_data_in[102]
port 55 nsew signal input
rlabel metal2 s 466550 0 466606 800 6 la_data_in[103]
port 56 nsew signal input
rlabel metal2 s 469862 0 469918 800 6 la_data_in[104]
port 57 nsew signal input
rlabel metal2 s 473174 0 473230 800 6 la_data_in[105]
port 58 nsew signal input
rlabel metal2 s 476486 0 476542 800 6 la_data_in[106]
port 59 nsew signal input
rlabel metal2 s 479798 0 479854 800 6 la_data_in[107]
port 60 nsew signal input
rlabel metal2 s 483110 0 483166 800 6 la_data_in[108]
port 61 nsew signal input
rlabel metal2 s 486422 0 486478 800 6 la_data_in[109]
port 62 nsew signal input
rlabel metal2 s 158534 0 158590 800 6 la_data_in[10]
port 63 nsew signal input
rlabel metal2 s 489734 0 489790 800 6 la_data_in[110]
port 64 nsew signal input
rlabel metal2 s 493046 0 493102 800 6 la_data_in[111]
port 65 nsew signal input
rlabel metal2 s 496358 0 496414 800 6 la_data_in[112]
port 66 nsew signal input
rlabel metal2 s 499670 0 499726 800 6 la_data_in[113]
port 67 nsew signal input
rlabel metal2 s 502982 0 503038 800 6 la_data_in[114]
port 68 nsew signal input
rlabel metal2 s 506294 0 506350 800 6 la_data_in[115]
port 69 nsew signal input
rlabel metal2 s 509606 0 509662 800 6 la_data_in[116]
port 70 nsew signal input
rlabel metal2 s 512918 0 512974 800 6 la_data_in[117]
port 71 nsew signal input
rlabel metal2 s 516230 0 516286 800 6 la_data_in[118]
port 72 nsew signal input
rlabel metal2 s 519542 0 519598 800 6 la_data_in[119]
port 73 nsew signal input
rlabel metal2 s 161846 0 161902 800 6 la_data_in[11]
port 74 nsew signal input
rlabel metal2 s 522854 0 522910 800 6 la_data_in[120]
port 75 nsew signal input
rlabel metal2 s 526166 0 526222 800 6 la_data_in[121]
port 76 nsew signal input
rlabel metal2 s 529478 0 529534 800 6 la_data_in[122]
port 77 nsew signal input
rlabel metal2 s 532790 0 532846 800 6 la_data_in[123]
port 78 nsew signal input
rlabel metal2 s 536102 0 536158 800 6 la_data_in[124]
port 79 nsew signal input
rlabel metal2 s 539414 0 539470 800 6 la_data_in[125]
port 80 nsew signal input
rlabel metal2 s 542726 0 542782 800 6 la_data_in[126]
port 81 nsew signal input
rlabel metal2 s 546038 0 546094 800 6 la_data_in[127]
port 82 nsew signal input
rlabel metal2 s 165158 0 165214 800 6 la_data_in[12]
port 83 nsew signal input
rlabel metal2 s 168470 0 168526 800 6 la_data_in[13]
port 84 nsew signal input
rlabel metal2 s 171782 0 171838 800 6 la_data_in[14]
port 85 nsew signal input
rlabel metal2 s 175094 0 175150 800 6 la_data_in[15]
port 86 nsew signal input
rlabel metal2 s 178406 0 178462 800 6 la_data_in[16]
port 87 nsew signal input
rlabel metal2 s 181718 0 181774 800 6 la_data_in[17]
port 88 nsew signal input
rlabel metal2 s 185030 0 185086 800 6 la_data_in[18]
port 89 nsew signal input
rlabel metal2 s 188342 0 188398 800 6 la_data_in[19]
port 90 nsew signal input
rlabel metal2 s 128726 0 128782 800 6 la_data_in[1]
port 91 nsew signal input
rlabel metal2 s 191654 0 191710 800 6 la_data_in[20]
port 92 nsew signal input
rlabel metal2 s 194966 0 195022 800 6 la_data_in[21]
port 93 nsew signal input
rlabel metal2 s 198278 0 198334 800 6 la_data_in[22]
port 94 nsew signal input
rlabel metal2 s 201590 0 201646 800 6 la_data_in[23]
port 95 nsew signal input
rlabel metal2 s 204902 0 204958 800 6 la_data_in[24]
port 96 nsew signal input
rlabel metal2 s 208214 0 208270 800 6 la_data_in[25]
port 97 nsew signal input
rlabel metal2 s 211526 0 211582 800 6 la_data_in[26]
port 98 nsew signal input
rlabel metal2 s 214838 0 214894 800 6 la_data_in[27]
port 99 nsew signal input
rlabel metal2 s 218150 0 218206 800 6 la_data_in[28]
port 100 nsew signal input
rlabel metal2 s 221462 0 221518 800 6 la_data_in[29]
port 101 nsew signal input
rlabel metal2 s 132038 0 132094 800 6 la_data_in[2]
port 102 nsew signal input
rlabel metal2 s 224774 0 224830 800 6 la_data_in[30]
port 103 nsew signal input
rlabel metal2 s 228086 0 228142 800 6 la_data_in[31]
port 104 nsew signal input
rlabel metal2 s 231398 0 231454 800 6 la_data_in[32]
port 105 nsew signal input
rlabel metal2 s 234710 0 234766 800 6 la_data_in[33]
port 106 nsew signal input
rlabel metal2 s 238022 0 238078 800 6 la_data_in[34]
port 107 nsew signal input
rlabel metal2 s 241334 0 241390 800 6 la_data_in[35]
port 108 nsew signal input
rlabel metal2 s 244646 0 244702 800 6 la_data_in[36]
port 109 nsew signal input
rlabel metal2 s 247958 0 248014 800 6 la_data_in[37]
port 110 nsew signal input
rlabel metal2 s 251270 0 251326 800 6 la_data_in[38]
port 111 nsew signal input
rlabel metal2 s 254582 0 254638 800 6 la_data_in[39]
port 112 nsew signal input
rlabel metal2 s 135350 0 135406 800 6 la_data_in[3]
port 113 nsew signal input
rlabel metal2 s 257894 0 257950 800 6 la_data_in[40]
port 114 nsew signal input
rlabel metal2 s 261206 0 261262 800 6 la_data_in[41]
port 115 nsew signal input
rlabel metal2 s 264518 0 264574 800 6 la_data_in[42]
port 116 nsew signal input
rlabel metal2 s 267830 0 267886 800 6 la_data_in[43]
port 117 nsew signal input
rlabel metal2 s 271142 0 271198 800 6 la_data_in[44]
port 118 nsew signal input
rlabel metal2 s 274454 0 274510 800 6 la_data_in[45]
port 119 nsew signal input
rlabel metal2 s 277766 0 277822 800 6 la_data_in[46]
port 120 nsew signal input
rlabel metal2 s 281078 0 281134 800 6 la_data_in[47]
port 121 nsew signal input
rlabel metal2 s 284390 0 284446 800 6 la_data_in[48]
port 122 nsew signal input
rlabel metal2 s 287702 0 287758 800 6 la_data_in[49]
port 123 nsew signal input
rlabel metal2 s 138662 0 138718 800 6 la_data_in[4]
port 124 nsew signal input
rlabel metal2 s 291014 0 291070 800 6 la_data_in[50]
port 125 nsew signal input
rlabel metal2 s 294326 0 294382 800 6 la_data_in[51]
port 126 nsew signal input
rlabel metal2 s 297638 0 297694 800 6 la_data_in[52]
port 127 nsew signal input
rlabel metal2 s 300950 0 301006 800 6 la_data_in[53]
port 128 nsew signal input
rlabel metal2 s 304262 0 304318 800 6 la_data_in[54]
port 129 nsew signal input
rlabel metal2 s 307574 0 307630 800 6 la_data_in[55]
port 130 nsew signal input
rlabel metal2 s 310886 0 310942 800 6 la_data_in[56]
port 131 nsew signal input
rlabel metal2 s 314198 0 314254 800 6 la_data_in[57]
port 132 nsew signal input
rlabel metal2 s 317510 0 317566 800 6 la_data_in[58]
port 133 nsew signal input
rlabel metal2 s 320822 0 320878 800 6 la_data_in[59]
port 134 nsew signal input
rlabel metal2 s 141974 0 142030 800 6 la_data_in[5]
port 135 nsew signal input
rlabel metal2 s 324134 0 324190 800 6 la_data_in[60]
port 136 nsew signal input
rlabel metal2 s 327446 0 327502 800 6 la_data_in[61]
port 137 nsew signal input
rlabel metal2 s 330758 0 330814 800 6 la_data_in[62]
port 138 nsew signal input
rlabel metal2 s 334070 0 334126 800 6 la_data_in[63]
port 139 nsew signal input
rlabel metal2 s 337382 0 337438 800 6 la_data_in[64]
port 140 nsew signal input
rlabel metal2 s 340694 0 340750 800 6 la_data_in[65]
port 141 nsew signal input
rlabel metal2 s 344006 0 344062 800 6 la_data_in[66]
port 142 nsew signal input
rlabel metal2 s 347318 0 347374 800 6 la_data_in[67]
port 143 nsew signal input
rlabel metal2 s 350630 0 350686 800 6 la_data_in[68]
port 144 nsew signal input
rlabel metal2 s 353942 0 353998 800 6 la_data_in[69]
port 145 nsew signal input
rlabel metal2 s 145286 0 145342 800 6 la_data_in[6]
port 146 nsew signal input
rlabel metal2 s 357254 0 357310 800 6 la_data_in[70]
port 147 nsew signal input
rlabel metal2 s 360566 0 360622 800 6 la_data_in[71]
port 148 nsew signal input
rlabel metal2 s 363878 0 363934 800 6 la_data_in[72]
port 149 nsew signal input
rlabel metal2 s 367190 0 367246 800 6 la_data_in[73]
port 150 nsew signal input
rlabel metal2 s 370502 0 370558 800 6 la_data_in[74]
port 151 nsew signal input
rlabel metal2 s 373814 0 373870 800 6 la_data_in[75]
port 152 nsew signal input
rlabel metal2 s 377126 0 377182 800 6 la_data_in[76]
port 153 nsew signal input
rlabel metal2 s 380438 0 380494 800 6 la_data_in[77]
port 154 nsew signal input
rlabel metal2 s 383750 0 383806 800 6 la_data_in[78]
port 155 nsew signal input
rlabel metal2 s 387062 0 387118 800 6 la_data_in[79]
port 156 nsew signal input
rlabel metal2 s 148598 0 148654 800 6 la_data_in[7]
port 157 nsew signal input
rlabel metal2 s 390374 0 390430 800 6 la_data_in[80]
port 158 nsew signal input
rlabel metal2 s 393686 0 393742 800 6 la_data_in[81]
port 159 nsew signal input
rlabel metal2 s 396998 0 397054 800 6 la_data_in[82]
port 160 nsew signal input
rlabel metal2 s 400310 0 400366 800 6 la_data_in[83]
port 161 nsew signal input
rlabel metal2 s 403622 0 403678 800 6 la_data_in[84]
port 162 nsew signal input
rlabel metal2 s 406934 0 406990 800 6 la_data_in[85]
port 163 nsew signal input
rlabel metal2 s 410246 0 410302 800 6 la_data_in[86]
port 164 nsew signal input
rlabel metal2 s 413558 0 413614 800 6 la_data_in[87]
port 165 nsew signal input
rlabel metal2 s 416870 0 416926 800 6 la_data_in[88]
port 166 nsew signal input
rlabel metal2 s 420182 0 420238 800 6 la_data_in[89]
port 167 nsew signal input
rlabel metal2 s 151910 0 151966 800 6 la_data_in[8]
port 168 nsew signal input
rlabel metal2 s 423494 0 423550 800 6 la_data_in[90]
port 169 nsew signal input
rlabel metal2 s 426806 0 426862 800 6 la_data_in[91]
port 170 nsew signal input
rlabel metal2 s 430118 0 430174 800 6 la_data_in[92]
port 171 nsew signal input
rlabel metal2 s 433430 0 433486 800 6 la_data_in[93]
port 172 nsew signal input
rlabel metal2 s 436742 0 436798 800 6 la_data_in[94]
port 173 nsew signal input
rlabel metal2 s 440054 0 440110 800 6 la_data_in[95]
port 174 nsew signal input
rlabel metal2 s 443366 0 443422 800 6 la_data_in[96]
port 175 nsew signal input
rlabel metal2 s 446678 0 446734 800 6 la_data_in[97]
port 176 nsew signal input
rlabel metal2 s 449990 0 450046 800 6 la_data_in[98]
port 177 nsew signal input
rlabel metal2 s 453302 0 453358 800 6 la_data_in[99]
port 178 nsew signal input
rlabel metal2 s 155222 0 155278 800 6 la_data_in[9]
port 179 nsew signal input
rlabel metal2 s 126518 0 126574 800 6 la_data_out[0]
port 180 nsew signal output
rlabel metal2 s 457718 0 457774 800 6 la_data_out[100]
port 181 nsew signal output
rlabel metal2 s 461030 0 461086 800 6 la_data_out[101]
port 182 nsew signal output
rlabel metal2 s 464342 0 464398 800 6 la_data_out[102]
port 183 nsew signal output
rlabel metal2 s 467654 0 467710 800 6 la_data_out[103]
port 184 nsew signal output
rlabel metal2 s 470966 0 471022 800 6 la_data_out[104]
port 185 nsew signal output
rlabel metal2 s 474278 0 474334 800 6 la_data_out[105]
port 186 nsew signal output
rlabel metal2 s 477590 0 477646 800 6 la_data_out[106]
port 187 nsew signal output
rlabel metal2 s 480902 0 480958 800 6 la_data_out[107]
port 188 nsew signal output
rlabel metal2 s 484214 0 484270 800 6 la_data_out[108]
port 189 nsew signal output
rlabel metal2 s 487526 0 487582 800 6 la_data_out[109]
port 190 nsew signal output
rlabel metal2 s 159638 0 159694 800 6 la_data_out[10]
port 191 nsew signal output
rlabel metal2 s 490838 0 490894 800 6 la_data_out[110]
port 192 nsew signal output
rlabel metal2 s 494150 0 494206 800 6 la_data_out[111]
port 193 nsew signal output
rlabel metal2 s 497462 0 497518 800 6 la_data_out[112]
port 194 nsew signal output
rlabel metal2 s 500774 0 500830 800 6 la_data_out[113]
port 195 nsew signal output
rlabel metal2 s 504086 0 504142 800 6 la_data_out[114]
port 196 nsew signal output
rlabel metal2 s 507398 0 507454 800 6 la_data_out[115]
port 197 nsew signal output
rlabel metal2 s 510710 0 510766 800 6 la_data_out[116]
port 198 nsew signal output
rlabel metal2 s 514022 0 514078 800 6 la_data_out[117]
port 199 nsew signal output
rlabel metal2 s 517334 0 517390 800 6 la_data_out[118]
port 200 nsew signal output
rlabel metal2 s 520646 0 520702 800 6 la_data_out[119]
port 201 nsew signal output
rlabel metal2 s 162950 0 163006 800 6 la_data_out[11]
port 202 nsew signal output
rlabel metal2 s 523958 0 524014 800 6 la_data_out[120]
port 203 nsew signal output
rlabel metal2 s 527270 0 527326 800 6 la_data_out[121]
port 204 nsew signal output
rlabel metal2 s 530582 0 530638 800 6 la_data_out[122]
port 205 nsew signal output
rlabel metal2 s 533894 0 533950 800 6 la_data_out[123]
port 206 nsew signal output
rlabel metal2 s 537206 0 537262 800 6 la_data_out[124]
port 207 nsew signal output
rlabel metal2 s 540518 0 540574 800 6 la_data_out[125]
port 208 nsew signal output
rlabel metal2 s 543830 0 543886 800 6 la_data_out[126]
port 209 nsew signal output
rlabel metal2 s 547142 0 547198 800 6 la_data_out[127]
port 210 nsew signal output
rlabel metal2 s 166262 0 166318 800 6 la_data_out[12]
port 211 nsew signal output
rlabel metal2 s 169574 0 169630 800 6 la_data_out[13]
port 212 nsew signal output
rlabel metal2 s 172886 0 172942 800 6 la_data_out[14]
port 213 nsew signal output
rlabel metal2 s 176198 0 176254 800 6 la_data_out[15]
port 214 nsew signal output
rlabel metal2 s 179510 0 179566 800 6 la_data_out[16]
port 215 nsew signal output
rlabel metal2 s 182822 0 182878 800 6 la_data_out[17]
port 216 nsew signal output
rlabel metal2 s 186134 0 186190 800 6 la_data_out[18]
port 217 nsew signal output
rlabel metal2 s 189446 0 189502 800 6 la_data_out[19]
port 218 nsew signal output
rlabel metal2 s 129830 0 129886 800 6 la_data_out[1]
port 219 nsew signal output
rlabel metal2 s 192758 0 192814 800 6 la_data_out[20]
port 220 nsew signal output
rlabel metal2 s 196070 0 196126 800 6 la_data_out[21]
port 221 nsew signal output
rlabel metal2 s 199382 0 199438 800 6 la_data_out[22]
port 222 nsew signal output
rlabel metal2 s 202694 0 202750 800 6 la_data_out[23]
port 223 nsew signal output
rlabel metal2 s 206006 0 206062 800 6 la_data_out[24]
port 224 nsew signal output
rlabel metal2 s 209318 0 209374 800 6 la_data_out[25]
port 225 nsew signal output
rlabel metal2 s 212630 0 212686 800 6 la_data_out[26]
port 226 nsew signal output
rlabel metal2 s 215942 0 215998 800 6 la_data_out[27]
port 227 nsew signal output
rlabel metal2 s 219254 0 219310 800 6 la_data_out[28]
port 228 nsew signal output
rlabel metal2 s 222566 0 222622 800 6 la_data_out[29]
port 229 nsew signal output
rlabel metal2 s 133142 0 133198 800 6 la_data_out[2]
port 230 nsew signal output
rlabel metal2 s 225878 0 225934 800 6 la_data_out[30]
port 231 nsew signal output
rlabel metal2 s 229190 0 229246 800 6 la_data_out[31]
port 232 nsew signal output
rlabel metal2 s 232502 0 232558 800 6 la_data_out[32]
port 233 nsew signal output
rlabel metal2 s 235814 0 235870 800 6 la_data_out[33]
port 234 nsew signal output
rlabel metal2 s 239126 0 239182 800 6 la_data_out[34]
port 235 nsew signal output
rlabel metal2 s 242438 0 242494 800 6 la_data_out[35]
port 236 nsew signal output
rlabel metal2 s 245750 0 245806 800 6 la_data_out[36]
port 237 nsew signal output
rlabel metal2 s 249062 0 249118 800 6 la_data_out[37]
port 238 nsew signal output
rlabel metal2 s 252374 0 252430 800 6 la_data_out[38]
port 239 nsew signal output
rlabel metal2 s 255686 0 255742 800 6 la_data_out[39]
port 240 nsew signal output
rlabel metal2 s 136454 0 136510 800 6 la_data_out[3]
port 241 nsew signal output
rlabel metal2 s 258998 0 259054 800 6 la_data_out[40]
port 242 nsew signal output
rlabel metal2 s 262310 0 262366 800 6 la_data_out[41]
port 243 nsew signal output
rlabel metal2 s 265622 0 265678 800 6 la_data_out[42]
port 244 nsew signal output
rlabel metal2 s 268934 0 268990 800 6 la_data_out[43]
port 245 nsew signal output
rlabel metal2 s 272246 0 272302 800 6 la_data_out[44]
port 246 nsew signal output
rlabel metal2 s 275558 0 275614 800 6 la_data_out[45]
port 247 nsew signal output
rlabel metal2 s 278870 0 278926 800 6 la_data_out[46]
port 248 nsew signal output
rlabel metal2 s 282182 0 282238 800 6 la_data_out[47]
port 249 nsew signal output
rlabel metal2 s 285494 0 285550 800 6 la_data_out[48]
port 250 nsew signal output
rlabel metal2 s 288806 0 288862 800 6 la_data_out[49]
port 251 nsew signal output
rlabel metal2 s 139766 0 139822 800 6 la_data_out[4]
port 252 nsew signal output
rlabel metal2 s 292118 0 292174 800 6 la_data_out[50]
port 253 nsew signal output
rlabel metal2 s 295430 0 295486 800 6 la_data_out[51]
port 254 nsew signal output
rlabel metal2 s 298742 0 298798 800 6 la_data_out[52]
port 255 nsew signal output
rlabel metal2 s 302054 0 302110 800 6 la_data_out[53]
port 256 nsew signal output
rlabel metal2 s 305366 0 305422 800 6 la_data_out[54]
port 257 nsew signal output
rlabel metal2 s 308678 0 308734 800 6 la_data_out[55]
port 258 nsew signal output
rlabel metal2 s 311990 0 312046 800 6 la_data_out[56]
port 259 nsew signal output
rlabel metal2 s 315302 0 315358 800 6 la_data_out[57]
port 260 nsew signal output
rlabel metal2 s 318614 0 318670 800 6 la_data_out[58]
port 261 nsew signal output
rlabel metal2 s 321926 0 321982 800 6 la_data_out[59]
port 262 nsew signal output
rlabel metal2 s 143078 0 143134 800 6 la_data_out[5]
port 263 nsew signal output
rlabel metal2 s 325238 0 325294 800 6 la_data_out[60]
port 264 nsew signal output
rlabel metal2 s 328550 0 328606 800 6 la_data_out[61]
port 265 nsew signal output
rlabel metal2 s 331862 0 331918 800 6 la_data_out[62]
port 266 nsew signal output
rlabel metal2 s 335174 0 335230 800 6 la_data_out[63]
port 267 nsew signal output
rlabel metal2 s 338486 0 338542 800 6 la_data_out[64]
port 268 nsew signal output
rlabel metal2 s 341798 0 341854 800 6 la_data_out[65]
port 269 nsew signal output
rlabel metal2 s 345110 0 345166 800 6 la_data_out[66]
port 270 nsew signal output
rlabel metal2 s 348422 0 348478 800 6 la_data_out[67]
port 271 nsew signal output
rlabel metal2 s 351734 0 351790 800 6 la_data_out[68]
port 272 nsew signal output
rlabel metal2 s 355046 0 355102 800 6 la_data_out[69]
port 273 nsew signal output
rlabel metal2 s 146390 0 146446 800 6 la_data_out[6]
port 274 nsew signal output
rlabel metal2 s 358358 0 358414 800 6 la_data_out[70]
port 275 nsew signal output
rlabel metal2 s 361670 0 361726 800 6 la_data_out[71]
port 276 nsew signal output
rlabel metal2 s 364982 0 365038 800 6 la_data_out[72]
port 277 nsew signal output
rlabel metal2 s 368294 0 368350 800 6 la_data_out[73]
port 278 nsew signal output
rlabel metal2 s 371606 0 371662 800 6 la_data_out[74]
port 279 nsew signal output
rlabel metal2 s 374918 0 374974 800 6 la_data_out[75]
port 280 nsew signal output
rlabel metal2 s 378230 0 378286 800 6 la_data_out[76]
port 281 nsew signal output
rlabel metal2 s 381542 0 381598 800 6 la_data_out[77]
port 282 nsew signal output
rlabel metal2 s 384854 0 384910 800 6 la_data_out[78]
port 283 nsew signal output
rlabel metal2 s 388166 0 388222 800 6 la_data_out[79]
port 284 nsew signal output
rlabel metal2 s 149702 0 149758 800 6 la_data_out[7]
port 285 nsew signal output
rlabel metal2 s 391478 0 391534 800 6 la_data_out[80]
port 286 nsew signal output
rlabel metal2 s 394790 0 394846 800 6 la_data_out[81]
port 287 nsew signal output
rlabel metal2 s 398102 0 398158 800 6 la_data_out[82]
port 288 nsew signal output
rlabel metal2 s 401414 0 401470 800 6 la_data_out[83]
port 289 nsew signal output
rlabel metal2 s 404726 0 404782 800 6 la_data_out[84]
port 290 nsew signal output
rlabel metal2 s 408038 0 408094 800 6 la_data_out[85]
port 291 nsew signal output
rlabel metal2 s 411350 0 411406 800 6 la_data_out[86]
port 292 nsew signal output
rlabel metal2 s 414662 0 414718 800 6 la_data_out[87]
port 293 nsew signal output
rlabel metal2 s 417974 0 418030 800 6 la_data_out[88]
port 294 nsew signal output
rlabel metal2 s 421286 0 421342 800 6 la_data_out[89]
port 295 nsew signal output
rlabel metal2 s 153014 0 153070 800 6 la_data_out[8]
port 296 nsew signal output
rlabel metal2 s 424598 0 424654 800 6 la_data_out[90]
port 297 nsew signal output
rlabel metal2 s 427910 0 427966 800 6 la_data_out[91]
port 298 nsew signal output
rlabel metal2 s 431222 0 431278 800 6 la_data_out[92]
port 299 nsew signal output
rlabel metal2 s 434534 0 434590 800 6 la_data_out[93]
port 300 nsew signal output
rlabel metal2 s 437846 0 437902 800 6 la_data_out[94]
port 301 nsew signal output
rlabel metal2 s 441158 0 441214 800 6 la_data_out[95]
port 302 nsew signal output
rlabel metal2 s 444470 0 444526 800 6 la_data_out[96]
port 303 nsew signal output
rlabel metal2 s 447782 0 447838 800 6 la_data_out[97]
port 304 nsew signal output
rlabel metal2 s 451094 0 451150 800 6 la_data_out[98]
port 305 nsew signal output
rlabel metal2 s 454406 0 454462 800 6 la_data_out[99]
port 306 nsew signal output
rlabel metal2 s 156326 0 156382 800 6 la_data_out[9]
port 307 nsew signal output
rlabel metal2 s 127622 0 127678 800 6 la_oenb[0]
port 308 nsew signal input
rlabel metal2 s 458822 0 458878 800 6 la_oenb[100]
port 309 nsew signal input
rlabel metal2 s 462134 0 462190 800 6 la_oenb[101]
port 310 nsew signal input
rlabel metal2 s 465446 0 465502 800 6 la_oenb[102]
port 311 nsew signal input
rlabel metal2 s 468758 0 468814 800 6 la_oenb[103]
port 312 nsew signal input
rlabel metal2 s 472070 0 472126 800 6 la_oenb[104]
port 313 nsew signal input
rlabel metal2 s 475382 0 475438 800 6 la_oenb[105]
port 314 nsew signal input
rlabel metal2 s 478694 0 478750 800 6 la_oenb[106]
port 315 nsew signal input
rlabel metal2 s 482006 0 482062 800 6 la_oenb[107]
port 316 nsew signal input
rlabel metal2 s 485318 0 485374 800 6 la_oenb[108]
port 317 nsew signal input
rlabel metal2 s 488630 0 488686 800 6 la_oenb[109]
port 318 nsew signal input
rlabel metal2 s 160742 0 160798 800 6 la_oenb[10]
port 319 nsew signal input
rlabel metal2 s 491942 0 491998 800 6 la_oenb[110]
port 320 nsew signal input
rlabel metal2 s 495254 0 495310 800 6 la_oenb[111]
port 321 nsew signal input
rlabel metal2 s 498566 0 498622 800 6 la_oenb[112]
port 322 nsew signal input
rlabel metal2 s 501878 0 501934 800 6 la_oenb[113]
port 323 nsew signal input
rlabel metal2 s 505190 0 505246 800 6 la_oenb[114]
port 324 nsew signal input
rlabel metal2 s 508502 0 508558 800 6 la_oenb[115]
port 325 nsew signal input
rlabel metal2 s 511814 0 511870 800 6 la_oenb[116]
port 326 nsew signal input
rlabel metal2 s 515126 0 515182 800 6 la_oenb[117]
port 327 nsew signal input
rlabel metal2 s 518438 0 518494 800 6 la_oenb[118]
port 328 nsew signal input
rlabel metal2 s 521750 0 521806 800 6 la_oenb[119]
port 329 nsew signal input
rlabel metal2 s 164054 0 164110 800 6 la_oenb[11]
port 330 nsew signal input
rlabel metal2 s 525062 0 525118 800 6 la_oenb[120]
port 331 nsew signal input
rlabel metal2 s 528374 0 528430 800 6 la_oenb[121]
port 332 nsew signal input
rlabel metal2 s 531686 0 531742 800 6 la_oenb[122]
port 333 nsew signal input
rlabel metal2 s 534998 0 535054 800 6 la_oenb[123]
port 334 nsew signal input
rlabel metal2 s 538310 0 538366 800 6 la_oenb[124]
port 335 nsew signal input
rlabel metal2 s 541622 0 541678 800 6 la_oenb[125]
port 336 nsew signal input
rlabel metal2 s 544934 0 544990 800 6 la_oenb[126]
port 337 nsew signal input
rlabel metal2 s 548246 0 548302 800 6 la_oenb[127]
port 338 nsew signal input
rlabel metal2 s 167366 0 167422 800 6 la_oenb[12]
port 339 nsew signal input
rlabel metal2 s 170678 0 170734 800 6 la_oenb[13]
port 340 nsew signal input
rlabel metal2 s 173990 0 174046 800 6 la_oenb[14]
port 341 nsew signal input
rlabel metal2 s 177302 0 177358 800 6 la_oenb[15]
port 342 nsew signal input
rlabel metal2 s 180614 0 180670 800 6 la_oenb[16]
port 343 nsew signal input
rlabel metal2 s 183926 0 183982 800 6 la_oenb[17]
port 344 nsew signal input
rlabel metal2 s 187238 0 187294 800 6 la_oenb[18]
port 345 nsew signal input
rlabel metal2 s 190550 0 190606 800 6 la_oenb[19]
port 346 nsew signal input
rlabel metal2 s 130934 0 130990 800 6 la_oenb[1]
port 347 nsew signal input
rlabel metal2 s 193862 0 193918 800 6 la_oenb[20]
port 348 nsew signal input
rlabel metal2 s 197174 0 197230 800 6 la_oenb[21]
port 349 nsew signal input
rlabel metal2 s 200486 0 200542 800 6 la_oenb[22]
port 350 nsew signal input
rlabel metal2 s 203798 0 203854 800 6 la_oenb[23]
port 351 nsew signal input
rlabel metal2 s 207110 0 207166 800 6 la_oenb[24]
port 352 nsew signal input
rlabel metal2 s 210422 0 210478 800 6 la_oenb[25]
port 353 nsew signal input
rlabel metal2 s 213734 0 213790 800 6 la_oenb[26]
port 354 nsew signal input
rlabel metal2 s 217046 0 217102 800 6 la_oenb[27]
port 355 nsew signal input
rlabel metal2 s 220358 0 220414 800 6 la_oenb[28]
port 356 nsew signal input
rlabel metal2 s 223670 0 223726 800 6 la_oenb[29]
port 357 nsew signal input
rlabel metal2 s 134246 0 134302 800 6 la_oenb[2]
port 358 nsew signal input
rlabel metal2 s 226982 0 227038 800 6 la_oenb[30]
port 359 nsew signal input
rlabel metal2 s 230294 0 230350 800 6 la_oenb[31]
port 360 nsew signal input
rlabel metal2 s 233606 0 233662 800 6 la_oenb[32]
port 361 nsew signal input
rlabel metal2 s 236918 0 236974 800 6 la_oenb[33]
port 362 nsew signal input
rlabel metal2 s 240230 0 240286 800 6 la_oenb[34]
port 363 nsew signal input
rlabel metal2 s 243542 0 243598 800 6 la_oenb[35]
port 364 nsew signal input
rlabel metal2 s 246854 0 246910 800 6 la_oenb[36]
port 365 nsew signal input
rlabel metal2 s 250166 0 250222 800 6 la_oenb[37]
port 366 nsew signal input
rlabel metal2 s 253478 0 253534 800 6 la_oenb[38]
port 367 nsew signal input
rlabel metal2 s 256790 0 256846 800 6 la_oenb[39]
port 368 nsew signal input
rlabel metal2 s 137558 0 137614 800 6 la_oenb[3]
port 369 nsew signal input
rlabel metal2 s 260102 0 260158 800 6 la_oenb[40]
port 370 nsew signal input
rlabel metal2 s 263414 0 263470 800 6 la_oenb[41]
port 371 nsew signal input
rlabel metal2 s 266726 0 266782 800 6 la_oenb[42]
port 372 nsew signal input
rlabel metal2 s 270038 0 270094 800 6 la_oenb[43]
port 373 nsew signal input
rlabel metal2 s 273350 0 273406 800 6 la_oenb[44]
port 374 nsew signal input
rlabel metal2 s 276662 0 276718 800 6 la_oenb[45]
port 375 nsew signal input
rlabel metal2 s 279974 0 280030 800 6 la_oenb[46]
port 376 nsew signal input
rlabel metal2 s 283286 0 283342 800 6 la_oenb[47]
port 377 nsew signal input
rlabel metal2 s 286598 0 286654 800 6 la_oenb[48]
port 378 nsew signal input
rlabel metal2 s 289910 0 289966 800 6 la_oenb[49]
port 379 nsew signal input
rlabel metal2 s 140870 0 140926 800 6 la_oenb[4]
port 380 nsew signal input
rlabel metal2 s 293222 0 293278 800 6 la_oenb[50]
port 381 nsew signal input
rlabel metal2 s 296534 0 296590 800 6 la_oenb[51]
port 382 nsew signal input
rlabel metal2 s 299846 0 299902 800 6 la_oenb[52]
port 383 nsew signal input
rlabel metal2 s 303158 0 303214 800 6 la_oenb[53]
port 384 nsew signal input
rlabel metal2 s 306470 0 306526 800 6 la_oenb[54]
port 385 nsew signal input
rlabel metal2 s 309782 0 309838 800 6 la_oenb[55]
port 386 nsew signal input
rlabel metal2 s 313094 0 313150 800 6 la_oenb[56]
port 387 nsew signal input
rlabel metal2 s 316406 0 316462 800 6 la_oenb[57]
port 388 nsew signal input
rlabel metal2 s 319718 0 319774 800 6 la_oenb[58]
port 389 nsew signal input
rlabel metal2 s 323030 0 323086 800 6 la_oenb[59]
port 390 nsew signal input
rlabel metal2 s 144182 0 144238 800 6 la_oenb[5]
port 391 nsew signal input
rlabel metal2 s 326342 0 326398 800 6 la_oenb[60]
port 392 nsew signal input
rlabel metal2 s 329654 0 329710 800 6 la_oenb[61]
port 393 nsew signal input
rlabel metal2 s 332966 0 333022 800 6 la_oenb[62]
port 394 nsew signal input
rlabel metal2 s 336278 0 336334 800 6 la_oenb[63]
port 395 nsew signal input
rlabel metal2 s 339590 0 339646 800 6 la_oenb[64]
port 396 nsew signal input
rlabel metal2 s 342902 0 342958 800 6 la_oenb[65]
port 397 nsew signal input
rlabel metal2 s 346214 0 346270 800 6 la_oenb[66]
port 398 nsew signal input
rlabel metal2 s 349526 0 349582 800 6 la_oenb[67]
port 399 nsew signal input
rlabel metal2 s 352838 0 352894 800 6 la_oenb[68]
port 400 nsew signal input
rlabel metal2 s 356150 0 356206 800 6 la_oenb[69]
port 401 nsew signal input
rlabel metal2 s 147494 0 147550 800 6 la_oenb[6]
port 402 nsew signal input
rlabel metal2 s 359462 0 359518 800 6 la_oenb[70]
port 403 nsew signal input
rlabel metal2 s 362774 0 362830 800 6 la_oenb[71]
port 404 nsew signal input
rlabel metal2 s 366086 0 366142 800 6 la_oenb[72]
port 405 nsew signal input
rlabel metal2 s 369398 0 369454 800 6 la_oenb[73]
port 406 nsew signal input
rlabel metal2 s 372710 0 372766 800 6 la_oenb[74]
port 407 nsew signal input
rlabel metal2 s 376022 0 376078 800 6 la_oenb[75]
port 408 nsew signal input
rlabel metal2 s 379334 0 379390 800 6 la_oenb[76]
port 409 nsew signal input
rlabel metal2 s 382646 0 382702 800 6 la_oenb[77]
port 410 nsew signal input
rlabel metal2 s 385958 0 386014 800 6 la_oenb[78]
port 411 nsew signal input
rlabel metal2 s 389270 0 389326 800 6 la_oenb[79]
port 412 nsew signal input
rlabel metal2 s 150806 0 150862 800 6 la_oenb[7]
port 413 nsew signal input
rlabel metal2 s 392582 0 392638 800 6 la_oenb[80]
port 414 nsew signal input
rlabel metal2 s 395894 0 395950 800 6 la_oenb[81]
port 415 nsew signal input
rlabel metal2 s 399206 0 399262 800 6 la_oenb[82]
port 416 nsew signal input
rlabel metal2 s 402518 0 402574 800 6 la_oenb[83]
port 417 nsew signal input
rlabel metal2 s 405830 0 405886 800 6 la_oenb[84]
port 418 nsew signal input
rlabel metal2 s 409142 0 409198 800 6 la_oenb[85]
port 419 nsew signal input
rlabel metal2 s 412454 0 412510 800 6 la_oenb[86]
port 420 nsew signal input
rlabel metal2 s 415766 0 415822 800 6 la_oenb[87]
port 421 nsew signal input
rlabel metal2 s 419078 0 419134 800 6 la_oenb[88]
port 422 nsew signal input
rlabel metal2 s 422390 0 422446 800 6 la_oenb[89]
port 423 nsew signal input
rlabel metal2 s 154118 0 154174 800 6 la_oenb[8]
port 424 nsew signal input
rlabel metal2 s 425702 0 425758 800 6 la_oenb[90]
port 425 nsew signal input
rlabel metal2 s 429014 0 429070 800 6 la_oenb[91]
port 426 nsew signal input
rlabel metal2 s 432326 0 432382 800 6 la_oenb[92]
port 427 nsew signal input
rlabel metal2 s 435638 0 435694 800 6 la_oenb[93]
port 428 nsew signal input
rlabel metal2 s 438950 0 439006 800 6 la_oenb[94]
port 429 nsew signal input
rlabel metal2 s 442262 0 442318 800 6 la_oenb[95]
port 430 nsew signal input
rlabel metal2 s 445574 0 445630 800 6 la_oenb[96]
port 431 nsew signal input
rlabel metal2 s 448886 0 448942 800 6 la_oenb[97]
port 432 nsew signal input
rlabel metal2 s 452198 0 452254 800 6 la_oenb[98]
port 433 nsew signal input
rlabel metal2 s 455510 0 455566 800 6 la_oenb[99]
port 434 nsew signal input
rlabel metal2 s 157430 0 157486 800 6 la_oenb[9]
port 435 nsew signal input
rlabel metal4 s 4208 2128 4528 349840 6 vccd1
port 436 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 349840 6 vccd1
port 436 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 349840 6 vccd1
port 436 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 349840 6 vccd1
port 436 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 349840 6 vccd1
port 436 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 349840 6 vccd1
port 436 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 349840 6 vccd1
port 436 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 349840 6 vccd1
port 436 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 349840 6 vccd1
port 436 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 349840 6 vccd1
port 436 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 349840 6 vccd1
port 436 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 349840 6 vccd1
port 436 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 349840 6 vccd1
port 436 nsew power bidirectional
rlabel metal4 s 403568 2128 403888 349840 6 vccd1
port 436 nsew power bidirectional
rlabel metal4 s 434288 2128 434608 349840 6 vccd1
port 436 nsew power bidirectional
rlabel metal4 s 465008 2128 465328 349840 6 vccd1
port 436 nsew power bidirectional
rlabel metal4 s 495728 2128 496048 349840 6 vccd1
port 436 nsew power bidirectional
rlabel metal4 s 526448 2128 526768 349840 6 vccd1
port 436 nsew power bidirectional
rlabel metal4 s 557168 2128 557488 349840 6 vccd1
port 436 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 349840 6 vssd1
port 437 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 349840 6 vssd1
port 437 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 349840 6 vssd1
port 437 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 349840 6 vssd1
port 437 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 349840 6 vssd1
port 437 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 349840 6 vssd1
port 437 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 349840 6 vssd1
port 437 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 349840 6 vssd1
port 437 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 349840 6 vssd1
port 437 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 349840 6 vssd1
port 437 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 349840 6 vssd1
port 437 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 349840 6 vssd1
port 437 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 349840 6 vssd1
port 437 nsew ground bidirectional
rlabel metal4 s 418928 2128 419248 349840 6 vssd1
port 437 nsew ground bidirectional
rlabel metal4 s 449648 2128 449968 349840 6 vssd1
port 437 nsew ground bidirectional
rlabel metal4 s 480368 2128 480688 349840 6 vssd1
port 437 nsew ground bidirectional
rlabel metal4 s 511088 2128 511408 349840 6 vssd1
port 437 nsew ground bidirectional
rlabel metal4 s 541808 2128 542128 349840 6 vssd1
port 437 nsew ground bidirectional
rlabel metal2 s 8390 0 8446 800 6 wb_clk_i
port 438 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 wb_rst_i
port 439 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 wbs_ack_o
port 440 nsew signal output
rlabel metal2 s 15014 0 15070 800 6 wbs_adr_i[0]
port 441 nsew signal input
rlabel metal2 s 52550 0 52606 800 6 wbs_adr_i[10]
port 442 nsew signal input
rlabel metal2 s 55862 0 55918 800 6 wbs_adr_i[11]
port 443 nsew signal input
rlabel metal2 s 59174 0 59230 800 6 wbs_adr_i[12]
port 444 nsew signal input
rlabel metal2 s 62486 0 62542 800 6 wbs_adr_i[13]
port 445 nsew signal input
rlabel metal2 s 65798 0 65854 800 6 wbs_adr_i[14]
port 446 nsew signal input
rlabel metal2 s 69110 0 69166 800 6 wbs_adr_i[15]
port 447 nsew signal input
rlabel metal2 s 72422 0 72478 800 6 wbs_adr_i[16]
port 448 nsew signal input
rlabel metal2 s 75734 0 75790 800 6 wbs_adr_i[17]
port 449 nsew signal input
rlabel metal2 s 79046 0 79102 800 6 wbs_adr_i[18]
port 450 nsew signal input
rlabel metal2 s 82358 0 82414 800 6 wbs_adr_i[19]
port 451 nsew signal input
rlabel metal2 s 19430 0 19486 800 6 wbs_adr_i[1]
port 452 nsew signal input
rlabel metal2 s 85670 0 85726 800 6 wbs_adr_i[20]
port 453 nsew signal input
rlabel metal2 s 88982 0 89038 800 6 wbs_adr_i[21]
port 454 nsew signal input
rlabel metal2 s 92294 0 92350 800 6 wbs_adr_i[22]
port 455 nsew signal input
rlabel metal2 s 95606 0 95662 800 6 wbs_adr_i[23]
port 456 nsew signal input
rlabel metal2 s 98918 0 98974 800 6 wbs_adr_i[24]
port 457 nsew signal input
rlabel metal2 s 102230 0 102286 800 6 wbs_adr_i[25]
port 458 nsew signal input
rlabel metal2 s 105542 0 105598 800 6 wbs_adr_i[26]
port 459 nsew signal input
rlabel metal2 s 108854 0 108910 800 6 wbs_adr_i[27]
port 460 nsew signal input
rlabel metal2 s 112166 0 112222 800 6 wbs_adr_i[28]
port 461 nsew signal input
rlabel metal2 s 115478 0 115534 800 6 wbs_adr_i[29]
port 462 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 wbs_adr_i[2]
port 463 nsew signal input
rlabel metal2 s 118790 0 118846 800 6 wbs_adr_i[30]
port 464 nsew signal input
rlabel metal2 s 122102 0 122158 800 6 wbs_adr_i[31]
port 465 nsew signal input
rlabel metal2 s 28262 0 28318 800 6 wbs_adr_i[3]
port 466 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 wbs_adr_i[4]
port 467 nsew signal input
rlabel metal2 s 35990 0 36046 800 6 wbs_adr_i[5]
port 468 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 wbs_adr_i[6]
port 469 nsew signal input
rlabel metal2 s 42614 0 42670 800 6 wbs_adr_i[7]
port 470 nsew signal input
rlabel metal2 s 45926 0 45982 800 6 wbs_adr_i[8]
port 471 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 wbs_adr_i[9]
port 472 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 wbs_cyc_i
port 473 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 wbs_dat_i[0]
port 474 nsew signal input
rlabel metal2 s 53654 0 53710 800 6 wbs_dat_i[10]
port 475 nsew signal input
rlabel metal2 s 56966 0 57022 800 6 wbs_dat_i[11]
port 476 nsew signal input
rlabel metal2 s 60278 0 60334 800 6 wbs_dat_i[12]
port 477 nsew signal input
rlabel metal2 s 63590 0 63646 800 6 wbs_dat_i[13]
port 478 nsew signal input
rlabel metal2 s 66902 0 66958 800 6 wbs_dat_i[14]
port 479 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 wbs_dat_i[15]
port 480 nsew signal input
rlabel metal2 s 73526 0 73582 800 6 wbs_dat_i[16]
port 481 nsew signal input
rlabel metal2 s 76838 0 76894 800 6 wbs_dat_i[17]
port 482 nsew signal input
rlabel metal2 s 80150 0 80206 800 6 wbs_dat_i[18]
port 483 nsew signal input
rlabel metal2 s 83462 0 83518 800 6 wbs_dat_i[19]
port 484 nsew signal input
rlabel metal2 s 20534 0 20590 800 6 wbs_dat_i[1]
port 485 nsew signal input
rlabel metal2 s 86774 0 86830 800 6 wbs_dat_i[20]
port 486 nsew signal input
rlabel metal2 s 90086 0 90142 800 6 wbs_dat_i[21]
port 487 nsew signal input
rlabel metal2 s 93398 0 93454 800 6 wbs_dat_i[22]
port 488 nsew signal input
rlabel metal2 s 96710 0 96766 800 6 wbs_dat_i[23]
port 489 nsew signal input
rlabel metal2 s 100022 0 100078 800 6 wbs_dat_i[24]
port 490 nsew signal input
rlabel metal2 s 103334 0 103390 800 6 wbs_dat_i[25]
port 491 nsew signal input
rlabel metal2 s 106646 0 106702 800 6 wbs_dat_i[26]
port 492 nsew signal input
rlabel metal2 s 109958 0 110014 800 6 wbs_dat_i[27]
port 493 nsew signal input
rlabel metal2 s 113270 0 113326 800 6 wbs_dat_i[28]
port 494 nsew signal input
rlabel metal2 s 116582 0 116638 800 6 wbs_dat_i[29]
port 495 nsew signal input
rlabel metal2 s 24950 0 25006 800 6 wbs_dat_i[2]
port 496 nsew signal input
rlabel metal2 s 119894 0 119950 800 6 wbs_dat_i[30]
port 497 nsew signal input
rlabel metal2 s 123206 0 123262 800 6 wbs_dat_i[31]
port 498 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 wbs_dat_i[3]
port 499 nsew signal input
rlabel metal2 s 33782 0 33838 800 6 wbs_dat_i[4]
port 500 nsew signal input
rlabel metal2 s 37094 0 37150 800 6 wbs_dat_i[5]
port 501 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 wbs_dat_i[6]
port 502 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 wbs_dat_i[7]
port 503 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 wbs_dat_i[8]
port 504 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 wbs_dat_i[9]
port 505 nsew signal input
rlabel metal2 s 17222 0 17278 800 6 wbs_dat_o[0]
port 506 nsew signal output
rlabel metal2 s 54758 0 54814 800 6 wbs_dat_o[10]
port 507 nsew signal output
rlabel metal2 s 58070 0 58126 800 6 wbs_dat_o[11]
port 508 nsew signal output
rlabel metal2 s 61382 0 61438 800 6 wbs_dat_o[12]
port 509 nsew signal output
rlabel metal2 s 64694 0 64750 800 6 wbs_dat_o[13]
port 510 nsew signal output
rlabel metal2 s 68006 0 68062 800 6 wbs_dat_o[14]
port 511 nsew signal output
rlabel metal2 s 71318 0 71374 800 6 wbs_dat_o[15]
port 512 nsew signal output
rlabel metal2 s 74630 0 74686 800 6 wbs_dat_o[16]
port 513 nsew signal output
rlabel metal2 s 77942 0 77998 800 6 wbs_dat_o[17]
port 514 nsew signal output
rlabel metal2 s 81254 0 81310 800 6 wbs_dat_o[18]
port 515 nsew signal output
rlabel metal2 s 84566 0 84622 800 6 wbs_dat_o[19]
port 516 nsew signal output
rlabel metal2 s 21638 0 21694 800 6 wbs_dat_o[1]
port 517 nsew signal output
rlabel metal2 s 87878 0 87934 800 6 wbs_dat_o[20]
port 518 nsew signal output
rlabel metal2 s 91190 0 91246 800 6 wbs_dat_o[21]
port 519 nsew signal output
rlabel metal2 s 94502 0 94558 800 6 wbs_dat_o[22]
port 520 nsew signal output
rlabel metal2 s 97814 0 97870 800 6 wbs_dat_o[23]
port 521 nsew signal output
rlabel metal2 s 101126 0 101182 800 6 wbs_dat_o[24]
port 522 nsew signal output
rlabel metal2 s 104438 0 104494 800 6 wbs_dat_o[25]
port 523 nsew signal output
rlabel metal2 s 107750 0 107806 800 6 wbs_dat_o[26]
port 524 nsew signal output
rlabel metal2 s 111062 0 111118 800 6 wbs_dat_o[27]
port 525 nsew signal output
rlabel metal2 s 114374 0 114430 800 6 wbs_dat_o[28]
port 526 nsew signal output
rlabel metal2 s 117686 0 117742 800 6 wbs_dat_o[29]
port 527 nsew signal output
rlabel metal2 s 26054 0 26110 800 6 wbs_dat_o[2]
port 528 nsew signal output
rlabel metal2 s 120998 0 121054 800 6 wbs_dat_o[30]
port 529 nsew signal output
rlabel metal2 s 124310 0 124366 800 6 wbs_dat_o[31]
port 530 nsew signal output
rlabel metal2 s 30470 0 30526 800 6 wbs_dat_o[3]
port 531 nsew signal output
rlabel metal2 s 34886 0 34942 800 6 wbs_dat_o[4]
port 532 nsew signal output
rlabel metal2 s 38198 0 38254 800 6 wbs_dat_o[5]
port 533 nsew signal output
rlabel metal2 s 41510 0 41566 800 6 wbs_dat_o[6]
port 534 nsew signal output
rlabel metal2 s 44822 0 44878 800 6 wbs_dat_o[7]
port 535 nsew signal output
rlabel metal2 s 48134 0 48190 800 6 wbs_dat_o[8]
port 536 nsew signal output
rlabel metal2 s 51446 0 51502 800 6 wbs_dat_o[9]
port 537 nsew signal output
rlabel metal2 s 18326 0 18382 800 6 wbs_sel_i[0]
port 538 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 wbs_sel_i[1]
port 539 nsew signal input
rlabel metal2 s 27158 0 27214 800 6 wbs_sel_i[2]
port 540 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 wbs_sel_i[3]
port 541 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 wbs_stb_i
port 542 nsew signal input
rlabel metal2 s 13910 0 13966 800 6 wbs_we_i
port 543 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 560000 352000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 53231150
string GDS_FILE /home/almund/git/c2s2/FFT_macro/openlane/user_proj_example/runs/23_05_01_18_26/results/signoff/user_proj_example.magic.gds
string GDS_START 389194
<< end >>

